// To be used inside controller.v

`define test 1'b0
`define test1 1'b1
