`include "defines.v"

module G1_Processor(
	input logic clk,
	input logic rst,
	input logic forward_EN
);
	
	logic writeEn, WB_EN_EXE, WB_EN_MEM, is_imm, ST, MEM_R_EN_EXE, hazard_detected, flagZ;
	logic brTaken, MEM_R_EN, MEM_W_EN, WB_EN;
	logic [`REG_FILE_ADDR_LEN-1:0] src1, src2, dest, dest_EXE, dest_MEM; 
	logic [`REG_FILE_SIZE-1:0]  writeVal, reg1, reg2, val1, val2;
	logic [`WORD_LEN-1:0] instruction_IF, instruction_ID; 
	logic [3:0] branch_comm;
	logic [`EXE_CMD_LEN-1:0] EXE_CMD;


	regFile rF(
		.clk(clk),
		.rst(rst),
		.writeEn(writeEn), //*
		.src1(src1),
		.src2(src2),
		.dest(dest),
		.writeVal(writeVal),
		
		.reg1(reg1),
		.reg2(reg2)
	);
	

	hazard_detection h_d(
		.src1_ID(src1),
		.src2_ID(src2),
		.dest_EXE(dest_EXE), //*
		.dest_MEM(dest_MEM), //*
		.op(instruction_ID[15:12]),
		.WB_EN_EXE(WB_EN_EXE), //*
		.WB_EN_MEM(WB_EN_MEM), //*
		.MEM_R_EN_EXE(MEM_R_EN_EXE), //*
		.forward_EN(forward_EN),
		.is_imm(is_imm),
		.ST(ST),
		
		
		.hazard_detected(hazard_detected)
	);
	

	IFStage ifS (
		.clk(clk),
		.rst(rst),
		.brTaken(brTaken),
		.brOffset(val2),
		.freeze(hazard_detected),
		.instruction(instruction_IF)
	);
	 
	 	
	IF_to_ID f2d(
		.clk(clk),
		.rst(rst),
		.flush(brTaken),
		.freeze(hazard_detected),
		.instructionIn(instruction_IF),
		.instruction(instruction_ID)
 	);
	

	ID id(
	  .hazard_detected(hazard_detected),
	  .flagZ(flagZ), //*
	  .instruction(instruction_ID), //*
	  .reg1(reg1),
	  .reg2(reg2),
	  
	  .brTaken(brTaken), 
	  .MEM_R_EN(MEM_R_EN), 
	  .MEM_W_EN(MEM_W_EN), 
	  .WB_EN(WB_EN), 
	  .is_imm_out(is_imm), 
	  .ST(ST), 
	  .EXE_CMD(EXE_CMD), 
	  .branch_comm(branch_comm), 
	  .src1(src1), 
	  .src2(src2), 
	  .val1(val1), 
	  .val2(val2)
  
  );


	logic alu_writeback_enable_out_pipe;
  logic alu_mem_read_enable_out_pipe;
  logic alu_mem_write_enable_out_pipe;
  logic [3:0] alu_instruction_dest_out_pipe;
  logic [23:0] alu_alu_result_out_pipe;
  logic [23:0] alu_write_data_out_pipe;
  ALU_to_MEM alu_to_mem(
    .rst(rst),
    .clk(clk),
    .writeback_enable(writeback_enable),
    .mem_read_enable(mem_read_enable),
    .mem_write_enable(mem_write_enable),
    .instruction_dest(instruction_dest),
    .alu_result(alu_result),
    .write_data(write_data),
    .writeback_enable_out(alu_writeback_enable_out_pipe),
    .mem_read_enable_out(alu_mem_read_enable_out_pipe),
    .mem_write_enable_out(alu_mem_write_enable_out_pipe),
    .instruction_dest_out(alu_instruction_dest_out_pipe),
    .alu_result_out(alu_alu_result_out_pipe),
    .write_data_out(alu_write_data_out_pipe)
  );


  logic memory_writeback_enable_out;
  logic memory_read_enable_out;
  logic [3:0] memory_instruction_dest_out;
  logic [23:0] memory_data_out;
  logic [23:0] memory_alu_result_out;
  logic [23:0] memory_data_b;
  memory_stage memory_stage(
    .rst(rst),
    .clk_a(clk),
    .clk_b(1'b0),
    .writeback_enable(alu_writeback_enable_out_pipe),
    .read_enable(alu_mem_read_enable_out_pipe),
    .write_enable(alu_mem_write_enable_out_pipe),
    .instruction_dest(alu_instruction_dest_out_pipe),
    .alu_result(alu_alu_result_out_pipe),
    .write_data_a(alu_write_data_out_pipe),
    .address_b(18'b0),
    .writeback_enable_out(memory_writeback_enable_out),
    .read_enable_out(memory_read_enable_out),
    .instruction_dest_out(memory_instruction_dest_out),
    .memory_out(memory_data_out),
    .alu_result_out(memory_alu_result_out),
    .read_data_b(memory_data_b)
  );


  logic memory_writeback_enable_out_pipe;
  logic memory_mem_read_enable_out_pipe;
  logic [3:0] memory_instruction_dest_out_pipe;
  logic [23:0] memory_mem_read_data_out_pipe;
  logic [23:0] memory_alu_result_pipe_out;
  MEM_to_WB mem_to_wb(
    .rst(rst),
    .clk(clk),
    .writeback_enable(memory_writeback_enable_out),
    .mem_read_enable(memory_read_enable_out),
    .instruction_dest(memory_instruction_dest_out),
    .mem_read_data(memory_data_out),
    .alu_result(memory_alu_result_out),
    .writeback_enable_out(memory_writeback_enable_out_pipe),
    .mem_read_enable_out(memory_mem_read_enable_out_pipe),
    .instruction_dest_out(memory_instruction_dest_out_pipe),
    .mem_read_data_out(memory_mem_read_data_out_pipe),
    .alu_result_out(memory_alu_result_pipe_out)
  );


  writeback_stage writeback_stage(
    .writeback_enable(memory_writeback_enable_out_pipe),
    .mem_read_enable(memory_mem_read_enable_out_pipe),
    .instruction_dest(memory_instruction_dest_out_pipe),
    .mem_read_data(memory_mem_read_data_out_pipe),
    .alu_result(memory_alu_result_pipe_out),
    .writeback_enable_out(writeEn),
    .instruction_dest_out(dest),
    .writeback_data_out(writeVal)
  );
endmodule 