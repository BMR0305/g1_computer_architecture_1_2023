module main(output logic a);
  assign a = 1;
endmodule